�� sr "it.polimi.is24am05.model.game.Gameޛmh�Q.9 I turnL 	gameStatet 0Lit/polimi/is24am05/model/enums/state/GameState;L goldDeckt $Lit/polimi/is24am05/model/deck/Deck;L playerst Ljava/util/List;L resourceDeckq ~ [ sharedObjectivest /[Lit/polimi/is24am05/model/objective/Objective;L winnersq ~ xp    ~r .it.polimi.is24am05.model.enums.state.GameState          xr java.lang.Enum          xpt GAMEsr "it.polimi.is24am05.model.deck.DeckP⁐��G L deckq ~ L visiblet Ljava/util/Set;xpsr java.util.LinkedList)S]J`�"  xpw   $~r /it.polimi.is24am05.model.card.goldCard.GoldCard          xq ~ t GC_046~q ~ t GC_076~q ~ t GC_061~q ~ t GC_044~q ~ t GC_065~q ~ t GC_080~q ~ t GC_063~q ~ t GC_067~q ~ t GC_054~q ~ t GC_071~q ~ t GC_048~q ~ t GC_066~q ~ t GC_059~q ~ t GC_058~q ~ t GC_074~q ~ t GC_070~q ~ t GC_064~q ~ t GC_057~q ~ t GC_060~q ~ t GC_078~q ~ t GC_069~q ~ t GC_056~q ~ t GC_055~q ~ t GC_073~q ~ t GC_062~q ~ t GC_079~q ~ t GC_051~q ~ t GC_068~q ~ t GC_043~q ~ t GC_052~q ~ t GC_049~q ~ t GC_072~q ~ t GC_047~q ~ t GC_041~q ~ t GC_045~q ~ t GC_050xsr java.util.HashSet�D�����4  xpw   ?@     ~q ~ t GC_077~q ~ t GC_053xsr java.util.ArrayListx����a� I sizexp   w   sr &it.polimi.is24am05.model.Player.Player�,V���| 
I pointsI satisfiedObjectiveCardsL colort &Lit/polimi/is24am05/model/enums/Color;L handq ~ L nicknamet Ljava/lang/String;L 	objectivet .Lit/polimi/is24am05/model/objective/Objective;[ objectivesHandq ~ L playAreat ,Lit/polimi/is24am05/model/playArea/PlayArea;L starterCardt 7Lit/polimi/is24am05/model/card/starterCard/StarterCard;L statet 2Lit/polimi/is24am05/model/enums/state/PlayerState;xp        ~r $it.polimi.is24am05.model.enums.Color          xq ~ t REDsq ~ ^   w   ~r 7it.polimi.is24am05.model.card.resourceCard.ResourceCard          xq ~ t RC_032~q ~ t GC_075~q ~ lt RC_018xt Leo~r ,it.polimi.is24am05.model.objective.Objective          xq ~ t O_101ur /[Lit.polimi.is24am05.model.objective.Objective;���_V�H  xp   q ~ u~q ~ tt O_087sr *it.polimi.is24am05.model.playArea.PlayAreaR����NN� 
I maxII maxJI minII minJI 	turnCountL blockedq ~ L frontierq ~ L orderedPlacementsq ~ L playAreat Ljava/util/Map;L visibleElementsq ~ |xp       ����       sq ~ Xw   ?@      xsq ~ Xw   ?@     sr 'it.polimi.is24am05.model.playArea.Tuple�<15�{�� I iI jxp��������sq ~ �      sq ~ �����    sq ~ �       sq ~ �����   sq ~ �   ����xsq ~ ^   w   sr -it.polimi.is24am05.model.card.side.PlacedSideb�ў�40 I 	turnCountL actualCoordt )Lit/polimi/is24am05/model/playArea/Tuple;L sidet )Lit/polimi/is24am05/model/card/side/Side;xp    sq ~ �        ~r 9it.polimi.is24am05.model.card.starterCard.StarterBackSide          xq ~ t SBS_085sq ~ �   sq ~ �����   ~r ;it.polimi.is24am05.model.card.resourceCard.ResourceBackSide          xq ~ t RBS_009xsr java.util.HashMap���`� F 
loadFactorI 	thresholdxp?@     w      q ~ �q ~ �q ~ �q ~ �xsq ~ �?@     w      ~r /it.polimi.is24am05.model.enums.element.Resource          xq ~ t FUNGIsr java.lang.Integer⠤���8 I valuexr java.lang.Number������  xp   ~q ~ �t ANIMALsq ~ �   ~r +it.polimi.is24am05.model.enums.element.Item          xq ~ t INKWELLsq ~ �    ~q ~ �t PLANTq ~ �~q ~ �t INSECTq ~ �~q ~ �t 
MANUSCRIPTq ~ �~q ~ �t QUILLq ~ �x~r 5it.polimi.is24am05.model.card.starterCard.StarterCard          xq ~ t SC_085~r 0it.polimi.is24am05.model.enums.state.PlayerState          xq ~ t PLACEsq ~ `       ~q ~ ht YELLOWsq ~ ^   w   ~q ~ lt RC_038~q ~ t GC_042~q ~ lt RC_030xt Andre~q ~ tt O_097uq ~ w   ~q ~ tt O_090q ~ �sq ~ {                 sq ~ Xw   ?@      xsq ~ Xw   ?@     sq ~ ���������sq ~ �      sq ~ �����   sq ~ �       sq ~ �   ����sq ~ �       xsq ~ ^   w   sq ~ �    sq ~ �        ~r :it.polimi.is24am05.model.card.starterCard.StarterFrontSide          xq ~ t SFS_083sq ~ �   sq ~ �      ~r <it.polimi.is24am05.model.card.resourceCard.ResourceFrontSide          xq ~ t RFS_020xsq ~ �?@     w      q ~ �q ~ �q ~ �q ~ �xsq ~ �?@     w      q ~ �q ~ �q ~ �q ~ �q ~ �q ~ �q ~ �sq ~ �   q ~ �q ~ �q ~ �q ~ �q ~ �q ~ �x~q ~ �t SC_083q ~ �xsq ~ 
sq ~ w    ~q ~ lt RC_003~q ~ lt RC_039~q ~ lt RC_005~q ~ lt RC_027~q ~ lt RC_034~q ~ lt RC_025~q ~ lt RC_007~q ~ lt RC_023~q ~ lt RC_010~q ~ lt RC_019~q ~ lt RC_026~q ~ lt RC_028~q ~ lt RC_013~q ~ lt RC_014~q ~ lt RC_001~q ~ lt RC_004~q ~ lt RC_006~q ~ lt RC_037~q ~ lt RC_031~q ~ lt RC_015~q ~ lt RC_021~q ~ lt RC_008~q ~ lt RC_011~q ~ lt RC_017~q ~ lt RC_033~q ~ lt RC_012~q ~ lt RC_024~q ~ lt RC_040~q ~ lt RC_022~q ~ lt RC_035~q ~ lt RC_029~q ~ lt RC_016xsq ~ Xw   ?@     ~q ~ lt RC_036~q ~ lt RC_002xuq ~ w   ~q ~ tt O_089~q ~ tt O_088sq ~ ^    w    x