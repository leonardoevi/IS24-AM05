�� sr "it.polimi.is24am05.model.game.GameM���( 	I turnL 	connectedt Ljava/util/Set;L 	gameStatet 0Lit/polimi/is24am05/model/enums/state/GameState;L goldDeckt $Lit/polimi/is24am05/model/deck/Deck;L lastGameStateq ~ L playerst Ljava/util/List;L resourceDeckq ~ [ sharedObjectivest /[Lit/polimi/is24am05/model/objective/Objective;L winnersq ~ xp    sr java.util.HashSet�D�����4  xpw   ?@     sr &it.polimi.is24am05.model.Player.Player�,V���| 
I pointsI satisfiedObjectiveCardsL colort &Lit/polimi/is24am05/model/enums/Color;L handq ~ L nicknamet Ljava/lang/String;L 	objectivet .Lit/polimi/is24am05/model/objective/Objective;[ objectivesHandq ~ L playAreat ,Lit/polimi/is24am05/model/playArea/PlayArea;L starterCardt 7Lit/polimi/is24am05/model/card/starterCard/StarterCard;L statet 2Lit/polimi/is24am05/model/enums/state/PlayerState;xp        ~r $it.polimi.is24am05.model.enums.Color          xr java.lang.Enum          xpt YELLOWsr java.util.ArrayListx����a� I sizexp   w   ~r 7it.polimi.is24am05.model.card.resourceCard.ResourceCard          xq ~ t RC_035~q ~ t RC_023~r /it.polimi.is24am05.model.card.goldCard.GoldCard          xq ~ t GC_065xt Leo~r ,it.polimi.is24am05.model.objective.Objective          xq ~ t O_095ur /[Lit.polimi.is24am05.model.objective.Objective;���_V�H  xp   ~q ~  t O_093q ~ !sr *it.polimi.is24am05.model.playArea.PlayAreaR����NN� 
I maxII maxJI minII minJI 	turnCountL blockedq ~ L frontierq ~ L orderedPlacementsq ~ L playAreat Ljava/util/Map;L visibleElementsq ~ (xp                   sq ~ w   ?@      xsq ~ w   ?@     sr 'it.polimi.is24am05.model.playArea.Tuple�<15�{�� I iI jxp��������sq ~ ,      sq ~ ,����   sq ~ ,   ����xsq ~    w   sr -it.polimi.is24am05.model.card.side.PlacedSideb�ў�40 I 	turnCountL actualCoordt )Lit/polimi/is24am05/model/playArea/Tuple;L sidet )Lit/polimi/is24am05/model/card/side/Side;xp    sq ~ ,        ~r :it.polimi.is24am05.model.card.starterCard.StarterFrontSide          xq ~ t SFS_082xsr java.util.HashMap���`� F 
loadFactorI 	thresholdxp?@     w      q ~ 6q ~ 5xsq ~ :?@     w      ~r /it.polimi.is24am05.model.enums.element.Resource          xq ~ t FUNGIsr java.lang.Integer⠤���8 I valuexr java.lang.Number������  xp   ~q ~ =t INSECTsq ~ @    ~r +it.polimi.is24am05.model.enums.element.Item          xq ~ t QUILLq ~ E~q ~ Ft 
MANUSCRIPTq ~ E~q ~ =t PLANTq ~ E~q ~ =t ANIMALsq ~ @   ~q ~ Ft INKWELLq ~ Ex~r 5it.polimi.is24am05.model.card.starterCard.StarterCard          xq ~ t SC_082~r 0it.polimi.is24am05.model.enums.state.PlayerState          xq ~ t PLACEsq ~ 	        ~q ~ t REDsq ~    w   ~q ~ t RC_012~q ~ t RC_005~q ~ t GC_056xt Andre~q ~  t O_102uq ~ #   q ~ c~q ~  t O_091sq ~ '                   sq ~ w   ?@      xsq ~ w   ?@     sq ~ ,��������sq ~ ,      sq ~ ,����   sq ~ ,   ����xsq ~    w   sq ~ 2    sq ~ ,        ~q ~ 7t SFS_084xsq ~ :?@     w      q ~ qq ~ pxsq ~ :?@     w      q ~ >q ~ Eq ~ Cq ~ Oq ~ Gq ~ Eq ~ Iq ~ Eq ~ Kq ~ Eq ~ Mq ~ Oq ~ Pq ~ Ex~q ~ Rt SC_084q ~ Vsq ~ 	        ~q ~ t GREENsq ~    w   ~q ~ t RC_030~q ~ t RC_013~q ~ t GC_049xt Manu~q ~  t O_099uq ~ #   q ~ �~q ~  t O_098sq ~ '                   sq ~ w   ?@     sq ~ ,      sq ~ ,   ����xsq ~ w   ?@     sq ~ ,��������sq ~ ,      sq ~ ,����   sq ~ ,   ����xsq ~    w   sq ~ 2    sq ~ ,        ~q ~ 7t SFS_085xsq ~ :?@     w      q ~ �q ~ �xsq ~ :?@     w      q ~ >q ~ Eq ~ Cq ~ Oq ~ Gq ~ Eq ~ Iq ~ Eq ~ Kq ~ Oq ~ Mq ~ Oq ~ Pq ~ Ex~q ~ Rt SC_085q ~ Vx~r .it.polimi.is24am05.model.enums.state.GameState          xq ~ t GAMEsr "it.polimi.is24am05.model.deck.DeckP⁐��G L deckq ~ L visibleq ~ xpsr java.util.LinkedList)S]J`�"  xpw   #~q ~ t GC_046~q ~ t GC_057~q ~ t GC_062~q ~ t GC_066~q ~ t GC_064~q ~ t GC_069~q ~ t GC_047~q ~ t GC_063~q ~ t GC_080~q ~ t GC_054~q ~ t GC_051~q ~ t GC_068~q ~ t GC_075~q ~ t GC_041~q ~ t GC_071~q ~ t GC_042~q ~ t GC_074~q ~ t GC_077~q ~ t GC_060~q ~ t GC_059~q ~ t GC_044~q ~ t GC_061~q ~ t GC_070~q ~ t GC_072~q ~ t GC_058~q ~ t GC_076~q ~ t GC_048~q ~ t GC_053~q ~ t GC_078~q ~ t GC_073~q ~ t GC_045~q ~ t GC_043~q ~ t GC_079~q ~ t GC_050~q ~ t GC_052xsq ~ w   ?@     ~q ~ t GC_067~q ~ t GC_055xpsq ~    w   q ~ Xq ~ xq ~ xsq ~ �sq ~ �w    ~q ~ t RC_017~q ~ t RC_038~q ~ t RC_022~q ~ t RC_031~q ~ t RC_036~q ~ t RC_018~q ~ t RC_021~q ~ t RC_034~q ~ t RC_029~q ~ t RC_014~q ~ t RC_026~q ~ t RC_024~q ~ t RC_032~q ~ t RC_040~q ~ t RC_007~q ~ t RC_037~q ~ t RC_019~q ~ t RC_020~q ~ t RC_033~q ~ t RC_003~q ~ t RC_039~q ~ t RC_016~q ~ t RC_009~q ~ t RC_001~q ~ t RC_004~q ~ t RC_025~q ~ t RC_002~q ~ t RC_027~q ~ t RC_006~q ~ t RC_011~q ~ t RC_028~q ~ t RC_015xsq ~ w   ?@     ~q ~ t RC_010~q ~ t RC_008xuq ~ #   ~q ~  t O_090~q ~  t O_096sq ~     w    x